library verilog;
use verilog.vl_types.all;
entity ComparadorMod7_vlg_vec_tst is
end ComparadorMod7_vlg_vec_tst;
