library verilog;
use verilog.vl_types.all;
entity circuitocombinacional_vlg_vec_tst is
end circuitocombinacional_vlg_vec_tst;
