library verilog;
use verilog.vl_types.all;
entity FFJK_vlg_vec_tst is
end FFJK_vlg_vec_tst;
