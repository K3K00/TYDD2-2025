library verilog;
use verilog.vl_types.all;
entity sumadorcompleto_vlg_vec_tst is
end sumadorcompleto_vlg_vec_tst;
