-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Thu Oct 23 14:38:41 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY esaeslacuestion IS 
	PORT
	(
		Hab_Dat :  IN  STD_LOGIC;
		SCL :  IN  STD_LOGIC;
		SDA :  IN  STD_LOGIC;
		fin_dato :  OUT  STD_LOGIC
	);
END esaeslacuestion;

ARCHITECTURE bdf_type OF esaeslacuestion IS 

COMPONENT contadormod7
	PORT(clock : IN STD_LOGIC;
		 cout : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT registro8bits
	PORT(clock : IN STD_LOGIC;
		 shiftin : IN STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_2 <= Hab_Dat AND SCL;


PORT MAP(clock => SYNTHESIZED_WIRE_2,
		 cout => fin_dato);


b2v_inst7 : registro8bits
PORT MAP(SDA => SDA,
		 shiftin => SYNTHESIZED_WIRE_2);


END bdf_type;