-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Sun Oct 19 12:04:49 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 
LIBRARY work;

ENTITY MultiplicadorSinSigno IS 
	PORT(	A0 :  IN  STD_LOGIC;
			A1 :  IN  STD_LOGIC;
			B0 :  IN  STD_LOGIC;
			B1 :  IN  STD_LOGIC;
			p0 :  OUT STD_LOGIC;
			p1 :  OUT STD_LOGIC;
			p2 :  OUT STD_LOGIC;
			p3 :  OUT STD_LOGIC
		);
END MultiplicadorSinSigno;

ARCHITECTURE bdf_type OF MultiplicadorSinSigno IS 

COMPONENT circuitocombinacional 
	PORT(a : IN STD_LOGIC;
		  b : IN STD_LOGIC;
		  cin : IN STD_LOGIC;
		  z : OUT STD_LOGIC;
		  cout : OUT STD_LOGIC
		  );
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC; --0V
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC; --0V
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_0 <= B0 AND A1;
SYNTHESIZED_WIRE_1 <= A0 AND B1;
SYNTHESIZED_WIRE_2 <= '0';
SYNTHESIZED_WIRE_4 <= A1 AND B1;
SYNTHESIZED_WIRE_5 <= '0';

p0 <= A0 AND B0;

b2v_inst2 : circuitocombinacional
PORT MAP(a => SYNTHESIZED_WIRE_0,
		   b => SYNTHESIZED_WIRE_1,
		   cin => SYNTHESIZED_WIRE_2,
		   z => p1,
		   cout => SYNTHESIZED_WIRE_3);

b2v_inst6 : circuitocombinacional
PORT MAP(a => SYNTHESIZED_WIRE_3,
		   b => SYNTHESIZED_WIRE_4,
		   cin => SYNTHESIZED_WIRE_5,
		   z => p2,
		   cout => p3);
END bdf_type;