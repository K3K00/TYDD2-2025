library verilog;
use verilog.vl_types.all;
entity esaeslacuestion_vlg_vec_tst is
end esaeslacuestion_vlg_vec_tst;
