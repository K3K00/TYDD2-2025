library verilog;
use verilog.vl_types.all;
entity MultiplicadorSinSigno_vlg_vec_tst is
end MultiplicadorSinSigno_vlg_vec_tst;
