-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Oct 21 16:37:48 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ImplementacionI2C IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clk : IN STD_LOGIC;
        SDA : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        Hab_Dir : OUT STD_LOGIC;
        Hab_Dat : OUT STD_LOGIC;
        ACK : OUT STD_LOGIC
    );
END ImplementacionI2C;

ARCHITECTURE BEHAVIOR OF ImplementacionI2C IS
    TYPE type_fstate IS (Oscioso,Guardadir,RyW,Acknowledge,Guardadato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clk,reg_fstate)
    BEGIN
        IF (clk='1' AND clk'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SDA,soy,fin_dir,fin_dato)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Oscioso;
            Hab_Dir <= '0';
            Hab_Dat <= '0';
            ACK <= '0';
        ELSE
            Hab_Dir <= '0';
            Hab_Dat <= '0';
            ACK <= '0';
            CASE fstate IS
                WHEN Oscioso =>
                    IF ((SDA = '1')) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((SDA = '0')) THEN
                        reg_fstate <= Guardadir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Oscioso;
                    END IF;

                    ACK <= '0';

                    Hab_Dir <= '0';

                    Hab_Dat <= '0';
                WHEN Guardadir =>
                    IF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= Oscioso;
                    ELSIF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= RyW;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= Guardadir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardadir;
                    END IF;

                    ACK <= '0';

                    Hab_Dir <= '1';

                    Hab_Dat <= '0';
                WHEN RyW =>
                    reg_fstate <= Acknowledge;

                    ACK <= '0';

                    Hab_Dir <= '0';

                    Hab_Dat <= '0';
                WHEN Acknowledge =>
                    reg_fstate <= Guardadato;

                    ACK <= '1';

                    Hab_Dir <= '0';

                    Hab_Dat <= '0';
                WHEN Guardadato =>
                    IF ((fin_dato = '1')) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((fin_dato = '0')) THEN
                        reg_fstate <= Guardadato;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardadato;
                    END IF;

                    ACK <= '0';

                    Hab_Dir <= '0';

                    Hab_Dat <= '1';
                WHEN OTHERS => 
                    Hab_Dir <= 'X';
                    Hab_Dat <= 'X';
                    ACK <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
