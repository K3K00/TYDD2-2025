library verilog;
use verilog.vl_types.all;
entity template_vlg_vec_tst is
end template_vlg_vec_tst;
