library verilog;
use verilog.vl_types.all;
entity sumadorcompleto_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end sumadorcompleto_vlg_check_tst;
