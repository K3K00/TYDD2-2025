library verilog;
use verilog.vl_types.all;
entity Template_vlg_check_tst is
    port(
        d_out           : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end Template_vlg_check_tst;
