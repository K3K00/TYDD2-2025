library verilog;
use verilog.vl_types.all;
entity FFJK_vlg_check_tst is
    port(
        Qout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FFJK_vlg_check_tst;
