library verilog;
use verilog.vl_types.all;
entity MultiplicadorSinSigno_vlg_check_tst is
    port(
        p0              : in     vl_logic;
        p1              : in     vl_logic;
        p2              : in     vl_logic;
        p3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MultiplicadorSinSigno_vlg_check_tst;
