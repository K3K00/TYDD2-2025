library verilog;
use verilog.vl_types.all;
entity seronoser_vlg_vec_tst is
end seronoser_vlg_vec_tst;
