library verilog;
use verilog.vl_types.all;
entity ImplementacionI2C_vlg_vec_tst is
end ImplementacionI2C_vlg_vec_tst;
