library verilog;
use verilog.vl_types.all;
entity esaeslacuestion_vlg_sample_tst is
    port(
        Hab_Dat         : in     vl_logic;
        SCL             : in     vl_logic;
        SDA             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end esaeslacuestion_vlg_sample_tst;
