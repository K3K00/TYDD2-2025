library verilog;
use verilog.vl_types.all;
entity esaeslacuestion_vlg_check_tst is
    port(
        fin_dato        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end esaeslacuestion_vlg_check_tst;
