library verilog;
use verilog.vl_types.all;
entity Esquematico_vlg_vec_tst is
end Esquematico_vlg_vec_tst;
