library verilog;
use verilog.vl_types.all;
entity MultiModyCA2_vlg_check_tst is
    port(
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        s2              : in     vl_logic;
        s3              : in     vl_logic;
        u0              : in     vl_logic;
        u1              : in     vl_logic;
        u2              : in     vl_logic;
        u3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MultiModyCA2_vlg_check_tst;
