library verilog;
use verilog.vl_types.all;
entity template_vlg_check_tst is
    port(
        dout            : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end template_vlg_check_tst;
