library verilog;
use verilog.vl_types.all;
entity StateTool_vlg_vec_tst is
end StateTool_vlg_vec_tst;
