library verilog;
use verilog.vl_types.all;
entity MultiModyCA2_vlg_vec_tst is
end MultiModyCA2_vlg_vec_tst;
