library verilog;
use verilog.vl_types.all;
entity MultiplicadorConSigno_vlg_vec_tst is
end MultiplicadorConSigno_vlg_vec_tst;
